`timescale 1ns / 1ps
module instruction_rom #( parameter WIDTH = 32)
(
	input logic CLK,
	input logic RESET,
	input logic [WIDTH-1:0] ADDRESS,
	output logic [WIDTH-1:0] INSTR
);

logic [WIDTH-1:0] temp_instr;

always@( posedge CLK or posedge RESET or posedge ADDRESS ) begin
	if( RESET ) temp_instr <= 32'bx;
	else begin
		case (ADDRESS/32'd4)
			32'd0: temp_instr <= 32'b11111100000000000000000000000000;
			32'd1: temp_instr <= 32'b00101100001010010100000000000000;
			32'd2: temp_instr <= 32'b00101100010010100100000000000000;
			32'd3: temp_instr <= 32'b11111100000000000000000000000000;
			32'd4: temp_instr <= 32'b11111100000000000000000000000000;
			32'd5: temp_instr <= 32'b11111100000000000000000000000000;
			32'd6: temp_instr <= 32'b11111100000000000000000000000000;
			32'd7: temp_instr <= 32'b11111100000000000000000000000000;
			32'd8: temp_instr <= 32'b00010000111000010001000000000001;
			32'd9: temp_instr <= 32'b11111100000000000000000000000000;
			32'd10: temp_instr <= 32'b11111100000000000000000000000000;
			32'd11: temp_instr <= 32'b11111100000000000000000000000000;
			32'd12: temp_instr <= 32'b11111100000000000000000000000000;
			32'd13: temp_instr <= 32'b11111100000000000000000000000000;
			32'd14: temp_instr <= 32'b00010001000001110001000000000001;
			32'd15: temp_instr <= 32'b11111100000000000000000000000000;
			32'd16: temp_instr <= 32'b11111100000000000000000000000000;
			32'd17: temp_instr <= 32'b11111100000000000000000000000000;
			32'd18: temp_instr <= 32'b11111100000000000000000000000000;
			32'd19: temp_instr <= 32'b11111100000000000000000000000000;
			default: temp_instr <= 32'b0;
		endcase
	end
end

assign INSTR = temp_instr;

endmodule